`include "riscv_opcodes.sv"

module riscv_alu
(
    input   [ 3:0] alu_op_i,
    input   [31:0] alu_a_i,
    input   [31:0] alu_b_i,
    output  [31:0] alu_c_o
);

begin

end
